
.param VDDVAL=3v

.global vdd vss gnd 

* supplies
vvdd vdd 0 dc VDDVAL
vgnd gnd 0 dc 0v
vss  vss 0 dc 0

.inc ./models

.subckt spi_blk in 
x1 in ctl nout nand
x2 nout mon inv
rctl ctl 0 1k 
rz z mon 10k
cz mon 0 4p
.ends

.subckt nand a b z
m3  z a c 0 n  l=0.3u w=3u as=1.0e-10 ad=1.0e-10 ps=0 pd=0
m4  c b  0  0 n  l=0.3u w=3u as=1.0e-10 ad=1.0e-10 ps=0 pd=0
m1  z b  vdd  vdd p l=0.5u w=5u as=1.0e-10 ad=1.0e-10 ps=0 pd=0
m2  z a  vdd  vdd p l=0.5u w=5u as=1.0e-10 ad=1.0e-10 ps=0 pd=0
.ends

.subckt inv a z 
m1 z a vdd vdd p l=0.5u w=5u as=1.0e-10 ad=1.0e-10 ps=0 pd=0  
m2 z a 0 0 n l=0.5u w=3u as=1.0e-10 ad=1.0e-10 ps=0 pd=0 
.ends
.print v(*)
.end
