bind fifo fifo_sva 
  #(.WIDTH(WIDTH),
    .DEPTH(DEPTH),
    .L2D(L2D))
i_fifo_bind
  (.*);
