bind fifo_ctrl fifo_ctrl_checker #(.DEPTH(DEPTH), .WIDTH(WIDTH)) chk(.*);
